// -----------------------------------------------------------------------------
// Left register for DES (32-bit by default)
// Next state during a round: L <= R_prev
// On init load:              L <= init_L (e.g., output of IP)
// -----------------------------------------------------------------------------

module left_reg #(
	parameter WIDTH = 32
)(
	input wire clk,
	input wire rst,
	input wire en,			// round enable (hold when 0)
	input wire load_init,		// load L_0 (initial value) when 1
	input wire [WIDTH-1:0] L_0,	// initial value
	input wire [WIDTH-1:0] R_prev,	// R_{n-1} (output of the previous round)
	output reg [WIDTH-1:0] L_curr	// current L
);

	wire [WIDTH-1:0] L_next = load_init ? L_0 :
				  en 	    ? R_prev :
					      L_curr;	// hold

	always @(posedge clk or negedge rst) begin
		if (!rst)
			L_curr <= {WIDTH{1'b0}};
		else
			L_curr <= L_next;
	end
endmodule
