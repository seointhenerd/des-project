// Module to perform S-box substitution (6 bits to 4 bits)

module SBox (
      input  wire [5:0] s_in,       // 6-bit input
      input  wire [2:0] box_num,    // S-box number (0-7)
      output reg  [3:0] s_out       // 4-bit output
);


 	// S-box 1
	/*localparam [3:0] S1 [0:63] = {
      	14, 4, 13, 1,  2, 15, 11, 8,  3, 10, 6, 12, 5,  9,  0, 7,
      	0, 15,  7, 4, 14,  2, 13, 1, 10,  6, 12, 11, 9,  5,  3, 8,
      	4,  1, 14, 8, 13,  6,  2, 11, 15, 12, 9,  7,  3, 10, 5, 0,
      	15, 12, 8, 2,  4,  9,  1,  7,  5, 11, 3, 14, 10, 0, 6, 13
	};

  	// S-box 2
  	localparam [3:0] S2 [0:63] = {
     	15,  1,  8, 14,  6, 11,  3,  4,  9,  7,  2, 13, 12,  0,  5, 10,
      	3, 13,  4,  7, 15,  2,  8, 14, 12,  0,  1, 10,  6,  9, 11,  5,
      	0, 14,  7, 11, 10,  4, 13,  1,  5,  8, 12,  6,  9,  3,  2, 15,
      	13,  8, 10,  1,  3, 15,  4,  2, 11,  6,  7, 12,  0,  5, 14,  9
  	};

  	// S-box 3
  	localparam [3:0] S3 [0:63] = {
      	10,  0,  9, 14,  6,  3, 15,  5,  1, 13, 12,  7, 11,  4,  2,  8,
      	13,  7,  0,  9,  3,  4,  6, 10,  2,  8,  5, 14, 12, 11, 15,  1,
      	13,  6,  4,  9,  8, 15,  3,  0, 11,  1,  2, 12,  5, 10, 14,  7,
      	1, 10, 13,  0,  6,  9,  8,  7,  4, 15, 14,  3, 11,  5,  2, 12
  	};

  	// S-box 4
  	localparam [3:0] S4 [0:63] = {
     	7, 13, 14,  3,  0,  6,  9, 10,  1,  2,  8,  5, 11, 12,  4, 15,
      	13,  8, 11,  5,  6, 15,  0,  3,  4,  7,  2, 12,  1, 10, 14,  9,
	10,  6,  9,  0, 12, 11,  7, 13, 15,  1,  3, 14,  5,  2,  8,  4,
      	3, 15,  0,  6, 10,  1, 13,  8,  9,  4,  5, 11, 12,  7,  2, 14
  	};

  	// S-box 5
  	localparam [3:0] S5 [0:63] = {
     	2, 12,  4,  1,  7, 10, 11,  6,  8,  5,  3, 15, 13,  0, 14,  9,
      	14, 11,  2, 12,  4,  7, 13,  1,  5,  0, 15, 10,  3,  9,  8,  6,
      	4,  2,  1, 11, 10, 13,  7,  8, 15,  9, 12,  5,  6,  3,  0, 14,
	11,  8, 12,  7,  1, 14,  2, 13,  6, 15,  0,  9, 10,  4,  5,  3
	};

  	// S-box 6
  	localparam [3:0] S6 [0:63] = {
      	12,  1, 10, 15,  9,  2,  6,  8,  0, 13,  3,  4, 14,  7,  5, 11,
      	10, 15,  4,  2,  7, 12,  9,  5,  6,  1, 13, 14,  0, 11,  3,  8,
      	9, 14, 15,  5,  2,  8, 12,  3,  7,  0,  4, 10,  1, 13, 11,  6,
	4,  3,  2, 12,  9,  5, 15, 10, 11, 14,  1,  7,  6,  0,  8, 13
  	};

  	// S-box 7
  	localparam [3:0] S7 [0:63] = {
      	4, 11,  2, 14, 15,  0,  8, 13,  3, 12,  9,  7,  5, 10,  6,  1,
      	13,  0, 11,  7,  4,  9,  1, 10, 14,  3,  5, 12,  2, 15,  8,  6,
      	1,  4, 11, 13, 12,  3,  7, 14, 10, 15,  6,  8,  0,  5,  9,  2,
      	6, 11, 13,  8,  1,  4, 10,  7,  9,  5,  0, 15, 14,  2,  3, 12
  	};

  	// S-box 8
  	localparam [3:0] S8 [0:63] = {
      	13,  2,  8,  4,  6, 15, 11,  1, 10,  9,  3, 14,  5,  0, 12,  7,
      	1, 15, 13,  8, 10,  3,  7,  4, 12,  5,  6, 11,  0, 14,  9,  2,
      	7, 11,  4,  1,  9, 12, 14,  2,  0,  6, 10, 13, 15,  3,  5,  8,
      	2,  1, 14,  7,  4, 10,  8, 13, 15, 12,  9,  0,  3,  5,  6, 11
  	};*/

	localparam [255:0] S1 = {
          4'd14, 4'd4, 4'd13, 4'd1,  4'd2, 4'd15, 4'd11, 4'd8,  4'd3, 4'd10, 4'd6, 4'd12, 4'd5,  4'd9,
  		4'd0, 4'd7,
          4'd0, 4'd15,  4'd7, 4'd4, 4'd14,  4'd2, 4'd13, 4'd1, 4'd10,  4'd6, 4'd12, 4'd11, 4'd9,  4'd5,
  		4'd3, 4'd8,
          4'd4,  4'd1, 4'd14, 4'd8, 4'd13,  4'd6,  4'd2, 4'd11, 4'd15, 4'd12, 4'd9,  4'd7,  4'd3, 4'd10,
  		4'd5, 4'd0,
          4'd15, 4'd12, 4'd8, 4'd2,  4'd4,  4'd9,  4'd1,  4'd7,  4'd5, 4'd11, 4'd3, 4'd14, 4'd10, 4'd0,
 		 4'd6, 4'd13
      };

	localparam [255:0] S2 = {
          4'd15,  4'd1,  4'd8, 4'd14,  4'd6, 4'd11,  4'd3,  4'd4,  4'd9,  4'd7,  4'd2, 4'd13, 4'd12,
  		4'd0,  4'd5, 4'd10,
          4'd3, 4'd13,  4'd4,  4'd7, 4'd15,  4'd2,  4'd8, 4'd14, 4'd12,  4'd0,  4'd1, 4'd10,  4'd6,  4'd9,
  		 4'd11,  4'd5,
          4'd0, 4'd14,  4'd7, 4'd11, 4'd10,  4'd4, 4'd13,  4'd1,  4'd5,  4'd8, 4'd12,  4'd6,  4'd9,  4'd3,
    		4'd2, 4'd15,
          4'd13,  4'd8, 4'd10,  4'd1,  4'd3, 4'd15,  4'd4,  4'd2, 4'd11,  4'd6,  4'd7, 4'd12,  4'd0,
  		4'd5, 4'd14,  4'd9
	};

	localparam [255:0] S3 = {
          4'd10,  4'd0,  4'd9, 4'd14,  4'd6,  4'd3, 4'd15,  4'd5,  4'd1, 4'd13, 4'd12,  4'd7, 4'd11,
  		4'd4,  4'd2,  4'd8,
          4'd13,  4'd7,  4'd0,  4'd9,  4'd3,  4'd4,  4'd6, 4'd10,  4'd2,  4'd8,  4'd5, 4'd14, 4'd12,
  		4'd11, 4'd15,  4'd1,
          4'd13,  4'd6,  4'd4,  4'd9,  4'd8, 4'd15,  4'd3,  4'd0, 4'd11,  4'd1,  4'd2, 4'd12,  4'd5,
  		4'd10, 4'd14,  4'd7,
          4'd1, 4'd10, 4'd13,  4'd0,  4'd6,  4'd9,  4'd8,  4'd7,  4'd4, 4'd15, 4'd14,  4'd3, 4'd11,  4'd5,
    		4'd2, 4'd12
	};

      localparam [255:0] S4 = {
          4'd7, 4'd13, 4'd14,  4'd3,  4'd0,  4'd6,  4'd9, 4'd10,  4'd1,  4'd2,  4'd8,  4'd5, 4'd11, 4'd12,
    4'd4, 4'd15,
          4'd13,  4'd8, 4'd11,  4'd5,  4'd6, 4'd15,  4'd0,  4'd3,  4'd4,  4'd7,  4'd2, 4'd12,  4'd1,
  4'd10, 4'd14,  4'd9,
          4'd10,  4'd6,  4'd9,  4'd0, 4'd12, 4'd11,  4'd7, 4'd13, 4'd15,  4'd1,  4'd3, 4'd14,  4'd5,
  4'd2,  4'd8,  4'd4,
          4'd3, 4'd15,  4'd0,  4'd6, 4'd10,  4'd1, 4'd13,  4'd8,  4'd9,  4'd4,  4'd5, 4'd11, 4'd12,  4'd7,
    4'd2, 4'd14
      };

      localparam [255:0] S5 = {
          4'd2, 4'd12,  4'd4,  4'd1,  4'd7, 4'd10, 4'd11,  4'd6,  4'd8,  4'd5,  4'd3, 4'd15, 4'd13,  4'd0,
   4'd14,  4'd9,
          4'd14, 4'd11,  4'd2, 4'd12,  4'd4,  4'd7, 4'd13,  4'd1,  4'd5,  4'd0, 4'd15, 4'd10,  4'd3,
  4'd9,  4'd8,  4'd6,
          4'd4,  4'd2,  4'd1, 4'd11, 4'd10, 4'd13,  4'd7,  4'd8, 4'd15,  4'd9, 4'd12,  4'd5,  4'd6,  4'd3,
    4'd0, 4'd14,
          4'd11,  4'd8, 4'd12,  4'd7,  4'd1, 4'd14,  4'd2, 4'd13,  4'd6, 4'd15,  4'd0,  4'd9, 4'd10,
  4'd4,  4'd5,  4'd3
      };

	localparam [255:0] S6 = {
          4'd12,  4'd1, 4'd10, 4'd15,  4'd9,  4'd2,  4'd6,  4'd8,  4'd0, 4'd13,  4'd3,  4'd4, 4'd14,
 		 4'd7,  4'd5, 4'd11,
          4'd10, 4'd15,  4'd4,  4'd2,  4'd7, 4'd12,  4'd9,  4'd5,  4'd6,  4'd1, 4'd13, 4'd14,  4'd0,
  		4'd11,  4'd3,  4'd8,
          4'd9, 4'd14, 4'd15,  4'd5,  4'd2,  4'd8, 4'd12,  4'd3,  4'd7,  4'd0,  4'd4, 4'd10,  4'd1, 4'd13,
   		4'd11,  4'd6,
          4'd4,  4'd3,  4'd2, 4'd12,  4'd9,  4'd5, 4'd15, 4'd10, 4'd11, 4'd14,  4'd1,  4'd7,  4'd6,  4'd0,
    		4'd8, 4'd13
	};

	localparam [255:0] S7 = {
          4'd4, 4'd11,  4'd2, 4'd14, 4'd15,  4'd0,  4'd8, 4'd13,  4'd3, 4'd12,  4'd9,  4'd7,  4'd5, 4'd10,
 		4'd6,  4'd1,
          4'd13,  4'd0, 4'd11,  4'd7,  4'd4,  4'd9,  4'd1, 4'd10, 4'd14,  4'd3,  4'd5, 4'd12,  4'd2,
  		4'd15,  4'd8,  4'd6,
          4'd1,  4'd4, 4'd11, 4'd13, 4'd12,  4'd3,  4'd7, 4'd14, 4'd10, 4'd15,  4'd6,  4'd8,  4'd0,  4'd5,
    		4'd9,  4'd2,
          4'd6, 4'd11, 4'd13,  4'd8,  4'd1,  4'd4, 4'd10,  4'd7,  4'd9,  4'd5,  4'd0, 4'd15, 4'd14,  4'd2,
    		4'd3, 4'd12
	};

	localparam [255:0] S8 = {
          4'd13,  4'd2,  4'd8,  4'd4,  4'd6, 4'd15, 4'd11,  4'd1, 4'd10,  4'd9,  4'd3, 4'd14,  4'd5,
  		4'd0, 4'd12,  4'd7,
          4'd1, 4'd15, 4'd13,  4'd8, 4'd10,  4'd3,  4'd7,  4'd4, 4'd12,  4'd5,  4'd6, 4'd11,  4'd0, 4'd14,
    		4'd9,  4'd2,
          4'd7, 4'd11,  4'd4,  4'd1,  4'd9, 4'd12, 4'd14,  4'd2,  4'd0,  4'd6, 4'd10, 4'd13, 4'd15,  4'd3,
    		4'd5,  4'd8,
          4'd2,  4'd1, 4'd14,  4'd7,  4'd4, 4'd10,  4'd8, 4'd13, 4'd15, 4'd12,  4'd9,  4'd0,  4'd3,  4'd5,
    		4'd6, 4'd11
	};


      wire [1:0] row;
      wire [3:0] col;
      wire [5:0] addr;

      assign row = {s_in[5], s_in[0]};
      assign col = s_in[4:1];
      assign addr = {row, col};

      // Select output using bit slicing
      always @(*) begin
          case (box_num)
              3'd0: s_out = S1[(63-addr)*4 +: 4];
              3'd1: s_out = S2[(63-addr)*4 +: 4];
              3'd2: s_out = S3[(63-addr)*4 +: 4];
              3'd3: s_out = S4[(63-addr)*4 +: 4];
              3'd4: s_out = S5[(63-addr)*4 +: 4];
              3'd5: s_out = S6[(63-addr)*4 +: 4];
              3'd6: s_out = S7[(63-addr)*4 +: 4];
              3'd7: s_out = S8[(63-addr)*4 +: 4];
              default: s_out = 4'd0;
          endcase
      end

  endmodule

