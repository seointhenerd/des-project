// Top-level Feistel function module. Implements f(R, K) = P(S(E(R) XOR K))

module Feistel_Function (
	input  wire [31:0] R_in,      // 32-bit right half
      	input  wire [47:0] subkey,    // 48-bit round subkey
     	output wire [31:0] f_out      // 32-bit output
);

     	wire [47:0] expansion_result; 
      	wire [47:0] xor_result;    
      	wire [31:0] sbox_result;  

      	// Stage 1: Expansion (32 bits to 48 bits)
      	Expansion exp_inst (
          .R_in(R_in),
          .E_out(expansion_result)
      	);

      	// Stage 2: XOR with subkey (48 bits)
      	assign xor_result = expansion_result ^ subkey;
	
      	// Stage 3: S-box substitution (48 bits to 32 bits)
      	SBoxArray sbox_inst (
          .xor_result(xor_result),
          .sbox_out(sbox_result)
      	);

      	// Stage 4: P-box permutation (32 bits to 32 bits)
      	PBox pbox_inst (
          .p_in(sbox_result),
          .p_out(f_out)
      	);

  endmodule
