`timescale 1ns / 1ps

module tb_Final_Permutation;

reg  [31:0] left_half;
reg  [31:0] right_half;
wire [63:0] output_text;

integer error_count;
reg [63:0] original_data;

Final_Permutation DUT (
    .left_half(left_half),
    .right_half(right_half),
    .output_text(output_text)
);


initial begin
    error_count = 0;

    // IP -> FP should be identity
    $display("Test: IP -> FP = identity check");
    original_data = 64'h0123_4567_89AB_CDEF;

    // Standard DES
    left_half  = 32'hCC00_CCFF;
    right_half = 32'hF0AA_F0AA;
    $display("left half: %h", left_half);
    $display("right half: %h", right_half);
    #10;

    if (output_text === original_data) begin
        $display("PASSED: FP(IP(x)) = x");
    end else begin
        $display("FAILED: FP is not inverse of IP");
        $display("  Expected: %h", original_data);
        $display("  Got:      %h", output_text);
        error_count = error_count + 1;
    end
    $display("");

    // Testing all zeros
    $display("Testing all zeros");
    left_half  = 32'h0000_0000;
    right_half = 32'h0000_0000;
    $display("left half: %h", left_half);
    $display("right half: %h", right_half);
    #10;

    if (output_text === 64'h0000_0000_0000_0000)
        $display("PASSED: All zeros");
    else begin
        $display("FAILED");
        error_count = error_count + 1;
    end
    $display("");

    // Testing all ones
    $display("Testing all ones");
    left_half  = 32'hFFFF_FFFF;
    right_half = 32'hFFFF_FFFF;
    $display("left half: %h", left_half);
    $display("right half: %h", right_half);
    #10;

    if (output_text === 64'hFFFF_FFFF_FFFF_FFFF)
        $display("PASSED: All ones");
    else begin
        $display("FAILED");
        error_count = error_count + 1;
    end
    $display("");


    // Testing known DES output
    $display("Testing known DES output");
    left_half  = 32'h4040_4040;
    right_half = 32'h0F0F_0F0F;
    #10;
    $display("Result = %h", output_text);
    $display("");

    // Testing Swap verification
    $display("Testing Swap verification");
    left_half  = 32'hAAAA_AAAA;
    right_half = 32'h5555_5555;
    #10;
    $display("Result = %h", output_text);
    $display("");

    $display("========================================");
    if (error_count == 0)
        $display("ALL TESTS PASSED!");
    else
        $display("%0d TEST(S) FAILED", error_count);
    $display("========================================\n");

    $finish;
end

endmodule
