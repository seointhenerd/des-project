module Control_State_Machine (
    input  wire clk,
    input  wire rst,
    input  wire start_encrypt,
    input  wire start_decrypt,
    input  wire [63:0] key,
    input  wire [63:0] input_text,
    
    output reg done_encrypt,
    output reg done_decrypt,
    output reg [63:0] output_text
);

    // State definitions
    localparam IDLE         = 3'b000;
    localparam INIT_PERM    = 3'b001;
    localparam ROUND_PROCESS = 3'b010;
    localparam FINAL_PERM   = 3'b011;
    localparam DONE         = 3'b100;
    
    reg [2:0] state;
    reg [3:0] round_counter;
    reg mode;  // 0=encrypt, 1=decrypt
    
    reg [31:0] left_reg, right_reg;
    reg [31:0] temp_reg;  // For swapping
    
    // Wires connecting to other modules
    wire [31:0] ip_left, ip_right;
    wire [63:0] fp_output;
    wire [31:0] f_output;
    
    // Subkey wires
    wire [47:0] k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, k16;
    
    // Current round subkey
    reg [47:0] current_subkey;
    
    // Initial Permutation
    Initial_Permutation ip_inst (
        .input_text(input_text),
        .left_half(ip_left),
        .right_half(ip_right)
    );
    
    // Subkey Generator
    key_schedule keygen_inst (
        .key(key),
        .k1(k1), .k2(k2), .k3(k3), .k4(k4),
        .k5(k5), .k6(k6), .k7(k7), .k8(k8),
        .k9(k9), .k10(k10), .k11(k11), .k12(k12),
        .k13(k13), .k14(k14), .k15(k15), .k16(k16)
    );
    
    // F-function
    Feistel_Function f_inst (
        .R_in(right_reg),
        .subkey(current_subkey),
        .f_out(f_output)
    );
    

    Final_Permutation fp_inst (
        .left_half(right_reg),
        .right_half(left_reg),
        .output_text(fp_output)
    );
    
    // Subkey selection - combinational
    always @(round_counter, mode, k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, k16) begin
        case (round_counter)
            4'd0:  current_subkey = mode ? k16 : k1;
            4'd1:  current_subkey = mode ? k15 : k2;
            4'd2:  current_subkey = mode ? k14 : k3;
            4'd3:  current_subkey = mode ? k13 : k4;
            4'd4:  current_subkey = mode ? k12 : k5;
            4'd5:  current_subkey = mode ? k11 : k6;
            4'd6:  current_subkey = mode ? k10 : k7;
            4'd7:  current_subkey = mode ? k9  : k8;
            4'd8:  current_subkey = mode ? k8  : k9;
            4'd9:  current_subkey = mode ? k7  : k10;
            4'd10: current_subkey = mode ? k6  : k11;
            4'd11: current_subkey = mode ? k5  : k12;
            4'd12: current_subkey = mode ? k4  : k13;
            4'd13: current_subkey = mode ? k3  : k14;
            4'd14: current_subkey = mode ? k2  : k15;
            4'd15: current_subkey = mode ? k1  : k16;
            default: current_subkey = k1;
        endcase
    end
    
    // FSM - sequential
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            state <= IDLE;
            round_counter <= 4'd0;
            done_encrypt <= 1'b0;
            done_decrypt <= 1'b0;
            left_reg <= 32'h0;
            right_reg <= 32'h0;
            output_text <= 64'h0;
            mode <= 1'b0;
        end else begin
            case (state)
                IDLE: begin
                    done_encrypt <= 1'b0;
                    done_decrypt <= 1'b0;
                    round_counter <= 4'd0;
                    
                    if (start_encrypt) begin
                        mode <= 1'b0;  // Encrypt
                        state <= INIT_PERM;
                    end else if (start_decrypt) begin
                        mode <= 1'b1;  // Decrypt
                        state <= INIT_PERM;
                    end
                end
                
                INIT_PERM: begin
                    // IP output -> registers
                    left_reg <= ip_left;
                    right_reg <= ip_right;
                    round_counter <= 4'd0;
                    state <= ROUND_PROCESS;
                end
                
                ROUND_PROCESS: begin
                    temp_reg <= right_reg;
                    left_reg <= right_reg;
                    right_reg <= left_reg ^ f_output;
                    
                    round_counter <= round_counter + 4'd1;
                    
                    // final permutation
                    if (round_counter == 4'd15) begin
                        state <= FINAL_PERM;
                    end
                end
                
                FINAL_PERM: begin
                    // FP output
                    output_text <= fp_output;
                    state <= DONE;
                end
                
                DONE: begin
                    if (mode == 1'b0) begin
                        done_encrypt <= 1'b1;
                    end else begin
                        done_decrypt <= 1'b1;
                    end
                    
                    if (!start_encrypt && !start_decrypt) begin
                        state <= IDLE;
                    end
                end
                
                default: state <= IDLE;
            endcase
        end
    end

endmodule